module x(input clk,a,b,output c); 

assign c = a & b & c;

endmodule